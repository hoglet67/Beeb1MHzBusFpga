library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity char_rom is
    generic (
        ADDR_WIDTH       : integer := 10;
        DATA_WIDTH       : integer := 8
    );
    port(
        clock    : in  std_logic;
        addressA : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
        QA       : out std_logic_vector(DATA_WIDTH-1 downto 0)
  );
end char_rom;

architecture RTL of char_rom is

    constant MEM_DEPTH : integer := 2**ADDR_WIDTH;

    type mem_type is array (0 to MEM_DEPTH-1) of unsigned(DATA_WIDTH-1 downto 0);

    shared variable mem : mem_type := (
        x"ff", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"ff", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"ff", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"ff", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"ff", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"ff", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"ff", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ff",
        x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80",
        x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40",
        x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20",
        x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10",
        x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08",
        x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04",
        x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02",
        x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"18", x"18", x"18", x"18", x"18", x"00", x"18", x"00",
        x"6c", x"6c", x"6c", x"00", x"00", x"00", x"00", x"00",
        x"36", x"36", x"7f", x"36", x"7f", x"36", x"36", x"00",
        x"0c", x"3f", x"68", x"3e", x"0b", x"7e", x"18", x"00",
        x"60", x"66", x"0c", x"18", x"30", x"66", x"06", x"00",
        x"38", x"6c", x"6c", x"38", x"6d", x"66", x"3b", x"00",
        x"0c", x"18", x"30", x"00", x"00", x"00", x"00", x"00",
        x"0c", x"18", x"30", x"30", x"30", x"18", x"0c", x"00",
        x"30", x"18", x"0c", x"0c", x"0c", x"18", x"30", x"00",
        x"00", x"18", x"7e", x"3c", x"7e", x"18", x"00", x"00",
        x"00", x"18", x"18", x"7e", x"18", x"18", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"30",
        x"00", x"00", x"00", x"7e", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00",
        x"00", x"06", x"0c", x"18", x"30", x"60", x"00", x"00",
        x"3c", x"66", x"6e", x"7e", x"76", x"66", x"3c", x"00",
        x"18", x"38", x"18", x"18", x"18", x"18", x"7e", x"00",
        x"3c", x"66", x"06", x"0c", x"18", x"30", x"7e", x"00",
        x"3c", x"66", x"06", x"1c", x"06", x"66", x"3c", x"00",
        x"0c", x"1c", x"3c", x"6c", x"7e", x"0c", x"0c", x"00",
        x"7e", x"60", x"7c", x"06", x"06", x"66", x"3c", x"00",
        x"1c", x"30", x"60", x"7c", x"66", x"66", x"3c", x"00",
        x"7e", x"06", x"0c", x"18", x"30", x"30", x"30", x"00",
        x"3c", x"66", x"66", x"3c", x"66", x"66", x"3c", x"00",
        x"3c", x"66", x"66", x"3e", x"06", x"0c", x"38", x"00",
        x"00", x"00", x"18", x"18", x"00", x"18", x"18", x"00",
        x"00", x"00", x"18", x"18", x"00", x"18", x"18", x"30",
        x"0c", x"18", x"30", x"60", x"30", x"18", x"0c", x"00",
        x"00", x"00", x"7e", x"00", x"7e", x"00", x"00", x"00",
        x"30", x"18", x"0c", x"06", x"0c", x"18", x"30", x"00",
        x"3c", x"66", x"0c", x"18", x"18", x"00", x"18", x"00",
        x"3c", x"66", x"6e", x"6a", x"6e", x"60", x"3c", x"00",
        x"3c", x"66", x"66", x"7e", x"66", x"66", x"66", x"00",
        x"7c", x"66", x"66", x"7c", x"66", x"66", x"7c", x"00",
        x"3c", x"66", x"60", x"60", x"60", x"66", x"3c", x"00",
        x"78", x"6c", x"66", x"66", x"66", x"6c", x"78", x"00",
        x"7e", x"60", x"60", x"7c", x"60", x"60", x"7e", x"00",
        x"7e", x"60", x"60", x"7c", x"60", x"60", x"60", x"00",
        x"3c", x"66", x"60", x"6e", x"66", x"66", x"3c", x"00",
        x"66", x"66", x"66", x"7e", x"66", x"66", x"66", x"00",
        x"7e", x"18", x"18", x"18", x"18", x"18", x"7e", x"00",
        x"3e", x"0c", x"0c", x"0c", x"0c", x"6c", x"38", x"00",
        x"66", x"6c", x"78", x"70", x"78", x"6c", x"66", x"00",
        x"60", x"60", x"60", x"60", x"60", x"60", x"7e", x"00",
        x"63", x"77", x"7f", x"6b", x"6b", x"63", x"63", x"00",
        x"66", x"66", x"76", x"7e", x"6e", x"66", x"66", x"00",
        x"3c", x"66", x"66", x"66", x"66", x"66", x"3c", x"00",
        x"7c", x"66", x"66", x"7c", x"60", x"60", x"60", x"00",
        x"3c", x"66", x"66", x"66", x"6a", x"6c", x"36", x"00",
        x"7c", x"66", x"66", x"7c", x"6c", x"66", x"66", x"00",
        x"3c", x"66", x"60", x"3c", x"06", x"66", x"3c", x"00",
        x"7e", x"18", x"18", x"18", x"18", x"18", x"18", x"00",
        x"66", x"66", x"66", x"66", x"66", x"66", x"3c", x"00",
        x"66", x"66", x"66", x"66", x"66", x"3c", x"18", x"00",
        x"63", x"63", x"6b", x"6b", x"7f", x"77", x"63", x"00",
        x"66", x"66", x"3c", x"18", x"3c", x"66", x"66", x"00",
        x"66", x"66", x"66", x"3c", x"18", x"18", x"18", x"00",
        x"7e", x"06", x"0c", x"18", x"30", x"60", x"7e", x"00",
        x"7c", x"60", x"60", x"60", x"60", x"60", x"7c", x"00",
        x"00", x"60", x"30", x"18", x"0c", x"06", x"00", x"00",
        x"3e", x"06", x"06", x"06", x"06", x"06", x"3e", x"00",
        x"18", x"3c", x"66", x"42", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"ff",
        x"1c", x"36", x"30", x"7c", x"30", x"30", x"7e", x"00",
        x"00", x"00", x"3c", x"06", x"3e", x"66", x"3e", x"00",
        x"60", x"60", x"7c", x"66", x"66", x"66", x"7c", x"00",
        x"00", x"00", x"3c", x"66", x"60", x"66", x"3c", x"00",
        x"06", x"06", x"3e", x"66", x"66", x"66", x"3e", x"00",
        x"00", x"00", x"3c", x"66", x"7e", x"60", x"3c", x"00",
        x"1c", x"30", x"30", x"7c", x"30", x"30", x"30", x"00",
        x"00", x"00", x"3e", x"66", x"66", x"3e", x"06", x"3c",
        x"60", x"60", x"7c", x"66", x"66", x"66", x"66", x"00",
        x"18", x"00", x"38", x"18", x"18", x"18", x"3c", x"00",
        x"18", x"00", x"38", x"18", x"18", x"18", x"18", x"70",
        x"60", x"60", x"66", x"6c", x"78", x"6c", x"66", x"00",
        x"38", x"18", x"18", x"18", x"18", x"18", x"3c", x"00",
        x"00", x"00", x"36", x"7f", x"6b", x"6b", x"63", x"00",
        x"00", x"00", x"7c", x"66", x"66", x"66", x"66", x"00",
        x"00", x"00", x"3c", x"66", x"66", x"66", x"3c", x"00",
        x"00", x"00", x"7c", x"66", x"66", x"7c", x"60", x"60",
        x"00", x"00", x"3e", x"66", x"66", x"3e", x"06", x"07",
        x"00", x"00", x"6c", x"76", x"60", x"60", x"60", x"00",
        x"00", x"00", x"3e", x"60", x"3c", x"06", x"7c", x"00",
        x"30", x"30", x"7c", x"30", x"30", x"30", x"1c", x"00",
        x"00", x"00", x"66", x"66", x"66", x"66", x"3e", x"00",
        x"00", x"00", x"66", x"66", x"66", x"3c", x"18", x"00",
        x"00", x"00", x"63", x"6b", x"6b", x"7f", x"36", x"00",
        x"00", x"00", x"66", x"3c", x"18", x"3c", x"66", x"00",
        x"00", x"00", x"66", x"66", x"66", x"3e", x"06", x"3c",
        x"00", x"00", x"7e", x"0c", x"18", x"30", x"7e", x"00",
        x"0c", x"18", x"18", x"70", x"18", x"18", x"0c", x"00",
        x"18", x"18", x"18", x"00", x"18", x"18", x"18", x"00",
        x"30", x"18", x"18", x"0e", x"18", x"18", x"30", x"00",
        x"31", x"6b", x"46", x"00", x"00", x"00", x"00", x"00",
        x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff", x"ff"
        );

begin

    process(clock) is
    begin
        if (rising_edge(clock)) then
            QA <= std_logic_vector(mem(to_integer(unsigned(addressA))));
        end if;
    end process;

end RTL;
